bind bool_proc bool_checker c0(.clk(clk), .rst(rst), .RT(RT), .RDY(RDY), .START(START), .ENDD(ENDD));
