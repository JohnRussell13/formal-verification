bind bool_proc bool_checker c0(.clk(clk), .rst(rst), .a(a), .y1(y1), .y2(y2), .z1(z1), .z2(z2));
