bind bool_proc bool_checker c0(.clk(clk), .rst(rst), .a(a), .b(b), .c(c), .d(d), .e(e), .f(f), .g(g), .h(h), .o1(o1), .o2(o2));
